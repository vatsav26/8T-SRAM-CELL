**8SRAM Read** 
* Power Supply 
Vdd 1 0 DC 1V         
* Control Signals 
Vwl 6 0 DC 0V        
Vbl 4 0 DC 0V         
Vblb 5 0 DC 0V       
Vrwl 7 0 PULSE(5 0 0 0 0 10u 20u)   
Vrbl 8 0 DC 1V        

* Models 
.model pmod pmos level=54 version=4.7 
.model nmod nmos level=54 version=4.7 

* Cross-coupled inverters (6T Core) 
M1 2 3 1 1 pmod W=20u L=1u     
M2 3 2 1 1 pmod W=20u L=1u    
M3 2 3 0 0 nmod W=10u L=1u     
M4 3 2 0 0 nmod W=10u L=1u    

* Write Access Transistors (disabled) 
M5 2 6 4 4 nmod W=10u L=1u     
M6 3 6 5 5 nmod W=10u L=1u     

* Read Access Transistors (enabled) 
M7 9 7 3 3 nmod W=10u L=1u     
M8 8 9 0 0 nmod W=10u L=1u     

* Simulation Control 
.control 
tran 1n 40u 
plot V(8) V(2) V(3)            
.endc 
.end
